`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:24:10 03/30/2016 
// Design Name: 
// Module Name:    Ext_32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Ext_32(
	input wire SEXT,
	input [15:0] imm_16,
	output [31:0] imm_32
	);

	assign imm_32 = SEXT==1 ? {{16{imm_16[15]}}, imm_16}:{16'h0, imm_16};
endmodule
