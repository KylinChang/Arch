`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:52:48 03/30/2016 
// Design Name: 
// Module Name:    IR_REG 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IR_REG(
input wire clk,
input wire rst,
input wire CE,
input wire[31:0] next_PC,
input wire[31:0] D,

output wire[31:0] IR_PC,
output reg[31:0] Q
    );


endmodule
