`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:37:39 04/17/2016 
// Design Name: 
// Module Name:    lui32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lui32(
input wire[31:0] imm,
output wire[31:0] o
    );

assign o[31:0] = imm[15:0];

endmodule
